// Signed integer division: result = signed(a) / signed(b)
module arith_divsi #(parameter int WIDTH = 32) (
    input  logic [WIDTH-1:0] a,
    input  logic [WIDTH-1:0] b,
    output logic [WIDTH-1:0] result
);
  assign result = $signed(a) / $signed(b);
endmodule
